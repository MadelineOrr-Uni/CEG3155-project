library ieee;
use ieee.std_logic_1164.all;

entity debugTLC is
	port (
	);
end entity;

architecture debugTLCArch of debugTLC is 

begin

end architecture;

